
`include "RegDef.vh"