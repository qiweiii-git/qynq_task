//*****************************************************************************
// RegDef.vh.
//
// Change History:
//  VER.   Author         DATE              Change Description
//  1.0    Qiwei Wu       Dec. 25, 2020     Initial Release
//*****************************************************************************

//*****************************************************************************
// reg defines
//*****************************************************************************
localparam FW_VER  = 0,
           LED_CTRL= 1,
           REG_CNT = 2;

//*****************************************************************************
// reg initialized value
//*****************************************************************************
wire [31:0] REG_INIT[0:REG_CNT-1];

assign REG_INIT[FW_VER]  = 32'h0006_0001;
assign REG_INIT[LED_CTRL] = 32'h0000_000F;
