
`include "RegDef.vh"
`include "QwiFmtDef.vh"